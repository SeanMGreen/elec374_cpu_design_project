module mem_data_reg (input [31:0] bus_mux_out,
                     input [31:0] m_data_in,
							input clr,
							input clk,
							input read,
							input mdrin,
							