module Datapath(input clock,
					 input r0out, r1out, r2out, r3out, r4out, r5out, r6out, r7out, r8out, 
                r9out, r10out, r11out, r12out, r13out, r14out, r15out, HIout, LOout,
					 Zhighout, Zlowout, PCout, MDRout, inportout, cout,
					 input [31:0] busmux_r0, busmux_r1, busmux_r2, busmux_r3, busmux_r4, 
					 busmux_r5, busmux_r6, busmux_r7, busmux_r8, busmux_r9, busmux_r10, 
					 busmux_r11, busmux_r12, busmux_r13, busmux_r14, busmux_r15, busmux_hi,
					 busmux_lo, busmux_zhigh, busmux_zlow, busmux_pc, busmux_mdr, busmux_inport, c_sign_extended);
					 

endmodule 
