module alu(a, b, alu_sel, c_hi, c_lo);
  input [31:0] a;
  input [31:0] b;
  input [3:0] alu_sel;
  output [31:0] c_hi;
  output [31:0] c_lo;
  wire c_in;
  wire c_out;
  wire [31:0] add_out;
  wire [31:0] sub_out;
  wire [63:0] mul_out;
  wire [63:0] div_out;
  wire [31:0] and_out;
  wire [31:0] or_out;
  wire [31:0] sr_out;
  wire [31:0] sl_out;
  wire [31:0] sra_out;
  wire [31:0] ror_out;
  wire [31:0] rol_out;
  wire [31:0] neg_out;
  wire [31:0] not_out;
  wire [30:0] mux0_temp2;
  wire [31:0] mux0_temp1;
  wire [31:0] mux0_temp0;
  wire [31:0] mux1_temp15;
  wire [31:0] mux1_temp14;
  wire [31:0] mux1_temp13;
  wire [31:0] mux1_temp12;
  wire [31:0] mux1_temp11;
  wire [31:0] mux1_temp10;
  wire [31:0] mux1_temp9;
  wire [31:0] mux1_temp8;
  wire [31:0] mux1_temp7;
  wire [31:0] mux1_temp4;
  wire [30:0] mux1_temp3;
  wire [31:0] mux1_temp2;
  wire [31:0] mux1_temp1;
  wire [31:0] mux1_temp0;
  wire enable;
  wire bo_in;
  wire bo_out;
  assign c_in = 0;
  assign mux0_temp2 = 0;
  assign mux0_temp1 = 0;
  assign mux0_temp0 = 0;
  assign mux1_temp15 = 0;
  assign mux1_temp14 = 0;
  assign mux1_temp13 = 0;
  assign mux1_temp12 = 0;
  assign mux1_temp11 = 0;
  assign mux1_temp10 = 0;
  assign mux1_temp9 = 0;
  assign mux1_temp8 = 0;
  assign mux1_temp7 = 0;
  assign mux1_temp4 = 0;
  assign mux1_temp3 = 0;
  assign mux1_temp2 = 0;
  assign mux1_temp1 = 0;
  assign mux1_temp0 = 0;
  assign bo_in = 1;
  rca_32_bit add(.c_out(c_out), .sum(add_out), .a(a), .b(b), .c_in(c_in));
  subtractor sub(.bo_out(bo_out), .d(sub_out), .a(a), .b(b), .bo_in(bo_in));
  booth_algorithm_32_bit mul(.m(a), .q(b), .p(mul_out));
  non_restoring_division  div(.q(a), .m(b), .output_val(div_out));
  AND_32_bit and_op(.a(a), .b(b), .c(and_out));
  OR_32_bit or_op(.a(a), .b(b), .c(or_out));
  shift_right(.a(a), .b(b), .c(sr_out));
  shift_left(.a(a), .b(b), .c(sl_out));
  shift_right_arithmetic(.a(a), .b(b), .c(sra_out));
  rotate_right(.a(a), .b(b), .c(ror_out));
  rotate_left(.a(a), .b(b), .c(rol_out));
  NEG_32_bit (.a(a), .b(neg_out));
  NOT_32_bit (.a(a), .b(not_out));
  mux16_to_1(.mux_out(c_lo), .data15(not_out), .data14(neg_out), .data13(rol_out), .data12(ror_out), .data11(shl_out), .data10(shra_out), .data9(shr_out), .data8(or_out), .data7(and_out), .data6(div_out[31:0]), .data5(mul_out[31:0]), .data4(sub_out), .data3(add_out), .data2(mux0_temp2), .data1(mux0_temp1), .data0(mux0_temp0));
  mux16_to_1(.mux_out(c_hi), .data15(mux1_temp15), .data14(mux1_temp14), .data13(mux1_temp13), .data12(mux1_temp12), .data11(mux1_temp11), .data10(mux1_temp10), .data9(mux1_temp9), .data8(mux1_temp8), .data7(mux1_temp7), .data6(div_out[63:32]), .data5(mul_out[63:32]), .data4(mux1_temp4), .data3({mux1_temp3, c_out}), .data2(mux1_temp2), .data1(mux1_temp1), .data0(mux1_temp0));
endmodule 
	
  
  
